library verilog;
use verilog.vl_types.all;
entity TrabalhoCircuitos_vlg_check_tst is
    port(
        SAIDA           : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end TrabalhoCircuitos_vlg_check_tst;
