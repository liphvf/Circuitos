library verilog;
use verilog.vl_types.all;
entity TrabalhoCircuitos_vlg_vec_tst is
end TrabalhoCircuitos_vlg_vec_tst;
